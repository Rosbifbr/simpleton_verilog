library verilog;
use verilog.vl_types.all;
entity simpleton_pitanga_vlg_vec_tst is
end simpleton_pitanga_vlg_vec_tst;
